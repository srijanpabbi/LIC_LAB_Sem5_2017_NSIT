*compensated non inverting amp
r1 0 2 1k
r2 2 3 1k
r4 3 4 1k
r3 6 4 1k 
x1 1 2 6 opamp1
x2 6 4 3 opamp1
*trans vin 1 0 sin(0 0.1 1k)
*ac
 vin 1 0 ac 0.1
*dc vin 1 0 dc 0
.lib C:\Users\LAB\Desktop\Srijan_ece3_2017\opamp1.lib
*.tran .9m 3m
*ac 
.ac dec 100 1 1000meg
*.dc vin -12 12 0.01
.probe
.end